`timescale 1ns / 1ps

//////////////////////////////////////////////////////////////////////////////////
//
// Created for Indiana University's E315 Class
//
// 
// Andrew Lukefahr
// lukefahr@iu.edu
//
// 2021-03-24
// 2020-04-27
//
//////////////////////////////////////////////////////////////////////////////////

module dot_20_10(

		// AXI4-Stream Interface
		input                           clk,
		input                           rst,

        // Incomming Matrix AXI4-Stream
		input [31:0]                    INPUT_AXIS_TDATA,
        input                           INPUT_AXIS_TLAST,
        input                           INPUT_AXIS_TVALID,
        output                          INPUT_AXIS_TREADY,
        
        // Outgoing Vector AXI4-Stream 		
		output [31:0]                   OUTPUT_AXIS_TDATA,
        output                          OUTPUT_AXIS_TLAST,
        output                          OUTPUT_AXIS_TVALID,
        input                           OUTPUT_AXIS_TREADY 

    );
    
// This is autogenerated. see python/dot_20_10.py for details. 
localparam ROWS = 20;
localparam COLS = 10;

localparam [31:0] weights [0:ROWS-1] [0:COLS-1] = '{
  '{
    $shortrealtobits(0.025832674),$shortrealtobits(0.031067913),$shortrealtobits(0.074954145),$shortrealtobits(0.069431275),
    $shortrealtobits(0.027941115),$shortrealtobits(-0.38890076),$shortrealtobits(0.033413205),$shortrealtobits(0.023418507),
    $shortrealtobits(0.06414384),$shortrealtobits(0.03908126)
  },
  '{
    $shortrealtobits(0.47429913),$shortrealtobits(-0.030727461),$shortrealtobits(-0.07559153),$shortrealtobits(-0.06562075),
    $shortrealtobits(-0.027017677),$shortrealtobits(-0.1192499),$shortrealtobits(-0.033655476),$shortrealtobits(-0.023151854),
    $shortrealtobits(-0.06256888),$shortrealtobits(-0.038519256)
  },
  '{
    $shortrealtobits(0.11026208),$shortrealtobits(-0.21939886),$shortrealtobits(0.13531552),$shortrealtobits(0.032739077),
    $shortrealtobits(-0.100836486),$shortrealtobits(0.0315356),$shortrealtobits(-0.070727594),$shortrealtobits(-0.060791247),
    $shortrealtobits(0.109173514),$shortrealtobits(-0.09761812)
  },
  '{
    $shortrealtobits(-0.09525199),$shortrealtobits(-0.015320993),$shortrealtobits(0.27705696),$shortrealtobits(0.29808667),
    $shortrealtobits(-0.0757019),$shortrealtobits(-0.35671774),$shortrealtobits(-0.36361465),$shortrealtobits(-0.19701016),
    $shortrealtobits(0.07038336),$shortrealtobits(-0.065721996)
  },
  '{
    $shortrealtobits(-0.0054014125),$shortrealtobits(-0.0017534702),$shortrealtobits(-0.02180146),$shortrealtobits(-0.043511778),
    $shortrealtobits(0.0126061505),$shortrealtobits(-0.06802737),$shortrealtobits(-0.022320164),$shortrealtobits(0.05773446),
    $shortrealtobits(0.0007781352),$shortrealtobits(0.093098156)
  },
  '{
    $shortrealtobits(0.15577213),$shortrealtobits(0.34477082),$shortrealtobits(0.090137675),$shortrealtobits(-0.31324303),
    $shortrealtobits(-0.3665532),$shortrealtobits(0.020112142),$shortrealtobits(-0.17536488),$shortrealtobits(0.30936924),
    $shortrealtobits(-0.33058545),$shortrealtobits(-0.14599612)
  },
  '{
    $shortrealtobits(0.0833357),$shortrealtobits(0.35463968),$shortrealtobits(0.034455944),$shortrealtobits(-0.17448412),
    $shortrealtobits(-0.14407434),$shortrealtobits(0.34011856),$shortrealtobits(-0.37385958),$shortrealtobits(0.21625571),
    $shortrealtobits(-0.31103995),$shortrealtobits(0.045323063)
  },
  '{
    $shortrealtobits(-0.02596514),$shortrealtobits(-0.034139764),$shortrealtobits(-0.074281424),$shortrealtobits(-0.06537479),
    $shortrealtobits(-0.027002666),$shortrealtobits(-0.12030753),$shortrealtobits(-0.032794163),$shortrealtobits(-0.022686793),
    $shortrealtobits(0.443038),$shortrealtobits(-0.04100036)
  },
  '{
    $shortrealtobits(-0.020247536),$shortrealtobits(-0.028367976),$shortrealtobits(-0.05547012),$shortrealtobits(-0.02299753),
    $shortrealtobits(0.4642982),$shortrealtobits(-0.049594223),$shortrealtobits(-0.012405541),$shortrealtobits(-0.08192114),
    $shortrealtobits(-0.063603744),$shortrealtobits(-0.13136235)
  },
  '{
    $shortrealtobits(-0.08965313),$shortrealtobits(-0.015638348),$shortrealtobits(0.31165576),$shortrealtobits(-0.0017556128),
    $shortrealtobits(0.22123784),$shortrealtobits(-0.29498687),$shortrealtobits(0.12892826),$shortrealtobits(-0.059905306),
    $shortrealtobits(-0.26068124),$shortrealtobits(-0.14420311)
  },
  '{
    $shortrealtobits(-0.021710042),$shortrealtobits(-0.029718418),$shortrealtobits(-0.05677786),$shortrealtobits(-0.024768198),
    $shortrealtobits(-0.037383515),$shortrealtobits(-0.052242942),$shortrealtobits(-0.0105619235),$shortrealtobits(0.42426327),
    $shortrealtobits(-0.062348627),$shortrealtobits(-0.12969314)
  },
  '{
    $shortrealtobits(-0.33830196),$shortrealtobits(-0.21303433),$shortrealtobits(-0.048951115),$shortrealtobits(0.25440967),
    $shortrealtobits(-0.22557631),$shortrealtobits(-0.09242142),$shortrealtobits(-0.055013154),$shortrealtobits(0.37846345),
    $shortrealtobits(0.2120045),$shortrealtobits(-0.2063289)
  },
  '{
    $shortrealtobits(-0.0014902132),$shortrealtobits(-0.5039727),$shortrealtobits(0.508414),$shortrealtobits(-0.001196809),
    $shortrealtobits(0.00043627736),$shortrealtobits(-0.0005926093),$shortrealtobits(-0.0012271563),$shortrealtobits(-0.00072608533),
    $shortrealtobits(-0.000416694),$shortrealtobits(2.0524347e-05)
  },
  '{
    $shortrealtobits(-0.026448617),$shortrealtobits(-0.031083299),$shortrealtobits(-0.07606366),$shortrealtobits(0.43673903),
    $shortrealtobits(-0.026514161),$shortrealtobits(-0.11752776),$shortrealtobits(-0.032170594),$shortrealtobits(-0.022210078),
    $shortrealtobits(-0.06506433),$shortrealtobits(-0.03911492)
  },
  '{
    $shortrealtobits(0.35377282),$shortrealtobits(-0.3778204),$shortrealtobits(0.29622322),$shortrealtobits(0.02397883),
    $shortrealtobits(-0.3820959),$shortrealtobits(-0.223997),$shortrealtobits(-0.16420537),$shortrealtobits(0.10098358),
    $shortrealtobits(-0.056816496),$shortrealtobits(-0.11162076)
  },
  '{
    $shortrealtobits(0.020578936),$shortrealtobits(0.028920183),$shortrealtobits(0.05403632),$shortrealtobits(0.023214692),
    $shortrealtobits(0.041436687),$shortrealtobits(0.049547866),$shortrealtobits(0.01047655),$shortrealtobits(0.0813296),
    $shortrealtobits(0.0643888),$shortrealtobits(-0.3736555)
  },
  '{
    $shortrealtobits(-0.02662784),$shortrealtobits(-0.03034657),$shortrealtobits(-0.0781744),$shortrealtobits(-0.06629315),
    $shortrealtobits(-0.027823025),$shortrealtobits(-0.11695455),$shortrealtobits(0.46898773),$shortrealtobits(-0.021602403),
    $shortrealtobits(-0.06392121),$shortrealtobits(-0.038148273)
  },
  '{
    $shortrealtobits(-0.21310297),$shortrealtobits(0.200328),$shortrealtobits(-0.2060856),$shortrealtobits(-0.25261205),
    $shortrealtobits(-0.13819245),$shortrealtobits(0.01940004),$shortrealtobits(0.019376138),$shortrealtobits(0.2770613),
    $shortrealtobits(-0.33503842),$shortrealtobits(-0.13916487)
  },
  '{
    $shortrealtobits(0.38198224),$shortrealtobits(-0.24366285),$shortrealtobits(0.120944664),$shortrealtobits(0.01898678),
    $shortrealtobits(0.20554696),$shortrealtobits(0.040481124),$shortrealtobits(0.23627168),$shortrealtobits(-0.28644764),
    $shortrealtobits(0.22857712),$shortrealtobits(0.4494442)
  },
  '{
    $shortrealtobits(-0.028221987),$shortrealtobits(-0.033350915),$shortrealtobits(0.43056083),$shortrealtobits(-0.06829891),
    $shortrealtobits(-0.02646765),$shortrealtobits(-0.117585674),$shortrealtobits(-0.03333983),$shortrealtobits(-0.022141851),
    $shortrealtobits(-0.06445468),$shortrealtobits(-0.037462544)
	}
};

    dot #(
        .ROWS(ROWS),
        .COLS(COLS)
    ) dot0 (
    
		// AXI4-Stream Interface
		.clk(clk),
		.rst(rst),
		
        .weights(weights),

        .INPUT_AXIS_TDATA(INPUT_AXIS_TDATA),
        .INPUT_AXIS_TLAST(INPUT_AXIS_TLAST),
        .INPUT_AXIS_TVALID(INPUT_AXIS_TVALID),
        .INPUT_AXIS_TREADY(INPUT_AXIS_TREADY),
                            
        .OUTPUT_AXIS_TDATA(OUTPUT_AXIS_TDATA),
        .OUTPUT_AXIS_TLAST(OUTPUT_AXIS_TLAST),
        .OUTPUT_AXIS_TVALID(OUTPUT_AXIS_TVALID),
        .OUTPUT_AXIS_TREADY(OUTPUT_AXIS_TREADY) 	

    );

    
endmodule
